VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dpll
  CLASS BLOCK ;
  FOREIGN dpll ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 596.000 225.310 600.000 ;
    END
  END clockp[1]
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 596.000 675.190 600.000 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 449.520 900.000 450.120 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END enable
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END resetb
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER nwell ;
        RECT 5.330 586.105 894.430 587.710 ;
        RECT 5.330 580.665 894.430 583.495 ;
        RECT 5.330 575.225 894.430 578.055 ;
        RECT 5.330 569.785 894.430 572.615 ;
        RECT 5.330 564.345 894.430 567.175 ;
        RECT 5.330 558.905 894.430 561.735 ;
        RECT 5.330 553.465 894.430 556.295 ;
        RECT 5.330 548.025 894.430 550.855 ;
        RECT 5.330 542.585 894.430 545.415 ;
        RECT 5.330 537.145 894.430 539.975 ;
        RECT 5.330 531.705 894.430 534.535 ;
        RECT 5.330 526.265 894.430 529.095 ;
        RECT 5.330 520.825 894.430 523.655 ;
        RECT 5.330 515.385 894.430 518.215 ;
        RECT 5.330 509.945 894.430 512.775 ;
        RECT 5.330 504.505 894.430 507.335 ;
        RECT 5.330 499.065 894.430 501.895 ;
        RECT 5.330 493.625 894.430 496.455 ;
        RECT 5.330 488.185 894.430 491.015 ;
        RECT 5.330 482.745 894.430 485.575 ;
        RECT 5.330 477.305 894.430 480.135 ;
        RECT 5.330 471.865 894.430 474.695 ;
        RECT 5.330 466.425 894.430 469.255 ;
        RECT 5.330 460.985 894.430 463.815 ;
        RECT 5.330 455.545 894.430 458.375 ;
        RECT 5.330 450.105 894.430 452.935 ;
        RECT 5.330 444.665 894.430 447.495 ;
        RECT 5.330 439.225 894.430 442.055 ;
        RECT 5.330 433.785 894.430 436.615 ;
        RECT 5.330 428.345 894.430 431.175 ;
        RECT 5.330 422.905 894.430 425.735 ;
        RECT 5.330 417.465 894.430 420.295 ;
        RECT 5.330 412.025 894.430 414.855 ;
        RECT 5.330 406.585 894.430 409.415 ;
        RECT 5.330 401.145 894.430 403.975 ;
        RECT 5.330 395.705 894.430 398.535 ;
        RECT 5.330 390.265 894.430 393.095 ;
        RECT 5.330 384.825 894.430 387.655 ;
        RECT 5.330 379.385 894.430 382.215 ;
        RECT 5.330 373.945 894.430 376.775 ;
        RECT 5.330 368.505 894.430 371.335 ;
        RECT 5.330 363.065 894.430 365.895 ;
        RECT 5.330 357.625 894.430 360.455 ;
        RECT 5.330 352.185 894.430 355.015 ;
        RECT 5.330 346.745 894.430 349.575 ;
        RECT 5.330 341.305 894.430 344.135 ;
        RECT 5.330 335.865 894.430 338.695 ;
        RECT 5.330 330.425 894.430 333.255 ;
        RECT 5.330 324.985 894.430 327.815 ;
        RECT 5.330 319.545 894.430 322.375 ;
        RECT 5.330 314.105 894.430 316.935 ;
        RECT 5.330 308.665 894.430 311.495 ;
        RECT 5.330 303.225 894.430 306.055 ;
        RECT 5.330 297.785 894.430 300.615 ;
        RECT 5.330 292.345 894.430 295.175 ;
        RECT 5.330 286.905 894.430 289.735 ;
        RECT 5.330 281.465 894.430 284.295 ;
        RECT 5.330 276.025 894.430 278.855 ;
        RECT 5.330 270.585 894.430 273.415 ;
        RECT 5.330 265.145 894.430 267.975 ;
        RECT 5.330 259.705 894.430 262.535 ;
        RECT 5.330 254.265 894.430 257.095 ;
        RECT 5.330 248.825 894.430 251.655 ;
        RECT 5.330 243.385 894.430 246.215 ;
        RECT 5.330 237.945 894.430 240.775 ;
        RECT 5.330 232.505 894.430 235.335 ;
        RECT 5.330 227.065 894.430 229.895 ;
        RECT 5.330 221.625 894.430 224.455 ;
        RECT 5.330 216.185 894.430 219.015 ;
        RECT 5.330 210.745 894.430 213.575 ;
        RECT 5.330 205.305 894.430 208.135 ;
        RECT 5.330 199.865 894.430 202.695 ;
        RECT 5.330 194.425 894.430 197.255 ;
        RECT 5.330 188.985 894.430 191.815 ;
        RECT 5.330 183.545 894.430 186.375 ;
        RECT 5.330 178.105 894.430 180.935 ;
        RECT 5.330 172.665 894.430 175.495 ;
        RECT 5.330 167.225 894.430 170.055 ;
        RECT 5.330 161.785 894.430 164.615 ;
        RECT 5.330 156.345 894.430 159.175 ;
        RECT 5.330 150.905 894.430 153.735 ;
        RECT 5.330 145.465 894.430 148.295 ;
        RECT 5.330 140.025 894.430 142.855 ;
        RECT 5.330 134.585 894.430 137.415 ;
        RECT 5.330 129.145 894.430 131.975 ;
        RECT 5.330 123.705 894.430 126.535 ;
        RECT 5.330 118.265 894.430 121.095 ;
        RECT 5.330 112.825 894.430 115.655 ;
        RECT 5.330 107.385 894.430 110.215 ;
        RECT 5.330 101.945 894.430 104.775 ;
        RECT 5.330 96.505 894.430 99.335 ;
        RECT 5.330 91.065 894.430 93.895 ;
        RECT 5.330 85.625 894.430 88.455 ;
        RECT 5.330 80.185 894.430 83.015 ;
        RECT 5.330 74.745 894.430 77.575 ;
        RECT 5.330 69.305 894.430 72.135 ;
        RECT 5.330 63.865 894.430 66.695 ;
        RECT 5.330 58.425 894.430 61.255 ;
        RECT 5.330 52.985 894.430 55.815 ;
        RECT 5.330 47.545 894.430 50.375 ;
        RECT 5.330 42.105 894.430 44.935 ;
        RECT 5.330 36.665 894.430 39.495 ;
        RECT 5.330 31.225 894.430 34.055 ;
        RECT 5.330 25.785 894.430 28.615 ;
        RECT 5.330 20.345 894.430 23.175 ;
        RECT 5.330 14.905 894.430 17.735 ;
        RECT 5.330 10.690 894.430 12.295 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 21.100 595.720 224.750 596.000 ;
        RECT 225.590 595.720 674.630 596.000 ;
        RECT 675.470 595.720 890.930 596.000 ;
        RECT 21.100 4.280 890.930 595.720 ;
        RECT 21.100 4.000 74.790 4.280 ;
        RECT 75.630 4.000 224.750 4.280 ;
        RECT 225.590 4.000 374.710 4.280 ;
        RECT 375.550 4.000 524.670 4.280 ;
        RECT 525.510 4.000 674.630 4.280 ;
        RECT 675.470 4.000 824.590 4.280 ;
        RECT 825.430 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 21.040 450.520 896.000 587.685 ;
        RECT 21.040 449.120 895.600 450.520 ;
        RECT 21.040 150.640 896.000 449.120 ;
        RECT 21.040 149.240 895.600 150.640 ;
        RECT 21.040 10.715 896.000 149.240 ;
      LAYER met4 ;
        RECT 523.775 140.255 541.585 167.785 ;
  END
END dpll
END LIBRARY

