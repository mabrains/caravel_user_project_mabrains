magic
tech sky130A
magscale 1 2
timestamp 1624041473
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 89994 119200 90050 120000
rect 22466 0 22522 800
rect 67454 0 67510 800
rect 112442 0 112498 800
rect 157430 0 157486 800
<< obsm2 >>
rect 1398 119144 89938 119200
rect 90106 119144 178092 119200
rect 1398 856 178092 119144
rect 1398 800 22410 856
rect 22578 800 67398 856
rect 67566 800 112386 856
rect 112554 800 157374 856
rect 157542 800 178092 856
<< metal3 >>
rect 179200 99968 180000 100088
rect 0 89904 800 90024
rect 179200 59984 180000 60104
rect 0 29928 800 30048
rect 179200 20000 180000 20120
<< obsm3 >>
rect 800 100168 179200 117537
rect 800 99888 179120 100168
rect 800 90104 179200 99888
rect 880 89824 179200 90104
rect 800 60184 179200 89824
rect 800 59904 179120 60184
rect 800 30128 179200 59904
rect 880 29848 179200 30128
rect 800 20200 179200 29848
rect 800 19920 179120 20200
rect 800 2143 179200 19920
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 95003 42739 96288 49197
rect 96768 42739 96948 49197
rect 97428 42739 97608 49197
rect 98088 42739 98268 49197
rect 98748 42739 99485 49197
<< labels >>
rlabel metal2 s 157430 0 157486 800 6 clockp[0]
port 1 nsew signal output
rlabel metal2 s 89994 119200 90050 120000 6 clockp[1]
port 2 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 div[0]
port 3 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 div[1]
port 4 nsew signal input
rlabel metal3 s 179200 20000 180000 20120 6 div[2]
port 5 nsew signal input
rlabel metal3 s 179200 59984 180000 60104 6 div[3]
port 6 nsew signal input
rlabel metal3 s 179200 99968 180000 100088 6 div[4]
port 7 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 enable
port 8 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 osc
port 9 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 resetb
port 10 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 11 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 17 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 20 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 21 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 23 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 24 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 25 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 26 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 27 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 28 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 29 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 30 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 31 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 32 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 33 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 34 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 35 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 36 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 37 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 38 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 39 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 40 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 41 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 42 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 43 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 44 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 45 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 46 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 47 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 48 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 49 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 50 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 51 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 52 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 53 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 54 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 55 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 56 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 57 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 58 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/dpll/runs/dpll/results/magic/dpll.gds
string GDS_END 5946434
string GDS_START 510002
<< end >>

